module hello_world;
  initial begin
    $display("Ciao CERN! Il simulatore funziona.");
    $finish;
  end
endmodule