// AUTOMATICALLY GENERATED - STABILIZED & CHECKED
// Format: Explicit Decimal (e.g. -8'd12)

// --- LAYER 1 ---
localparam signed [7:0] L1_N1_W1 = 8'd127;
localparam signed [7:0] L1_N1_W2 = 8'd127;
localparam signed [7:0] L1_N1_B  = -8'd128;
localparam signed [7:0] L1_N2_W1 = 8'd0;
localparam signed [7:0] L1_N2_W2 = 8'd0;
localparam signed [7:0] L1_N2_B  = -8'd128;
localparam signed [7:0] L1_N3_W1 = -8'd128;
localparam signed [7:0] L1_N3_W2 = -8'd128;
localparam signed [7:0] L1_N3_B  = 8'd127;

// --- LAYER 2 ---
localparam signed [7:0] L2_W1 = 8'd127;
localparam signed [7:0] L2_W2 = 8'd0;
localparam signed [7:0] L2_W3 = -8'd128;
localparam signed [7:0] L2_B  = -8'd14;
