`timescale 1ns / 1ps

module layer_1 (
    input clk,
    input rst,
    input signed [7:0] input_energy,
    input signed [7:0] input_isol,
    output signed [15:0] n1_out,
    output signed [15:0] n2_out,
    output signed [15:0] n3_out
);

    // --- SIDELOADING INTELLIGENCE ---
    // This command tells Verilog: "Stop guessing and read the Python script."
    // It pulls in the 'localparam' definitions generated by master_config.py
    `include "weights.vh"

    // --- PATCHING THE MATRIX (Mapping Params to Wires) ---
    
    // NEURON 1: The First Responder
    wire signed [7:0] w1_1 = L1_N1_W1; // Downloaded from weights.vh
    wire signed [7:0] w1_2 = L1_N1_W2;
    wire signed [7:0] b1   = L1_N1_B;

    // NEURON 2: The Skeptic
    wire signed [7:0] w2_1 = L1_N2_W1;
    wire signed [7:0] w2_2 = L1_N2_W2;
    wire signed [7:0] b2   = L1_N2_B;

    // NEURON 3: The Wildcard
    wire signed [7:0] w3_1 = L1_N3_W1;
    wire signed [7:0] w3_2 = L1_N3_W2;
    wire signed [7:0] b3   = L1_N3_B;

    // --- THE ENGINE ROOM (3 Neurons in a trenchcoat) ---
    neuron N1 (.clk(clk), .rst(rst), .x1(input_energy), .x2(input_isol), .w1(w1_1), .w2(w1_2), .b(b1), .y(n1_out));
    neuron N2 (.clk(clk), .rst(rst), .x1(input_energy), .x2(input_isol), .w1(w2_1), .w2(w2_2), .b(b2), .y(n2_out));
    neuron N3 (.clk(clk), .rst(rst), .x1(input_energy), .x2(input_isol), .w1(w3_1), .w2(w3_2), .b(b3), .y(n3_out));

endmodule