`timescale 1ns / 1ps

module layer_2 (
    input signed [15:0] n1,     // Input from Neuron 1: The Optimist
    input signed [15:0] n2,     // Input from Neuron 2: The Pessimist
    input signed [15:0] n3,     // Input from Neuron 3: The Wildcard
    output reg trigger,         // The Verdict: 1 = NOBEL PRIZE, 0 = TRASH
    output reg signed [31:0] score // The raw confidence score (for debugging insecurities)
);

    // --- IMPORTING THE HIVE MIND ---
    // This command opens the portal to the Python dimension.
    // It loads the magic numbers generated by master_config.py
    `include "weights.vh"

    // --- MAPPING THE DNA TO THE BODY ---
    // Extracting the specific genes (parameters) for this layer.
    wire signed [7:0] w1 = L2_W1;
    wire signed [7:0] w2 = L2_W2;
    wire signed [7:0] w3 = L2_W3;
    wire signed [7:0] b  = L2_B;

    always @(*) begin
        // --- THE JUDGMENT DAY ---
        // Summing up the opinions of the previous layer.
        // We use 32 bits because overflow is for amateurs.
        score = (n1 * w1) + (n2 * w2) + (n3 * w3) + b;

        // --- THE DECISION ---
        // If the score is positive, we found the Higgs. 
        // If negative, it's just cosmic background static.
        if (score > 0) 
            trigger = 1'b1; // FIRE! (Call Stockholm)
        else 
            trigger = 1'b0; // Silence. (Move along, nothing to see here)
    end

endmodule